package test_parameters_pkg;

    // typedef enums

    // parameters


endpackage