// Any further package imports:
import macro_pkg::*;

interface dp_sink_if(clk);
    string name_1, name_2, name_3;

    // modport DUT (
    //     input ctl
    // );
endinterface
