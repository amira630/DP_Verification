package dp_tl_agent_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Includes:
    `include "dp_source_config.svh"
    `include "dp_tl_sequencer.svh"
    `include "dp_tl_driver.svh"
    `include "dp_tl_monitor.svh"
    `include "dp_tl_agent.svh"

endpackage
