package dp_tl_agent_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Any further package imports:
    import dp_transactions_pkg::*;
    import test_parameters_pkg::*;
    
    // Includes:
    `include "dp_tl_sequencer.svh"
    `include "dp_tl_driver.svh"
    `include "dp_tl_monitor.svh"
    `include "dp_tl_agent.svh"

endpackage
