package dp_transactions_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import test_parameters_pkg::*;
    
    // Includes:
    `include "dp_source_config.svh"
    `include "dp_tl_sequence_item.svh"
    `include "dp_sink_sequence_item.svh"
    `include "dp_ref_transaction.svh"

endpackage