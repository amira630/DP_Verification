interface dp_sink_if(input clk);
    string name_1, name_2, name_3;

    // modport DUT (
    //     input ctl
    // );
endinterface
