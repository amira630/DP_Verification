interface DP_SINK_if(clk);
    // ... rest of the code
endinterface