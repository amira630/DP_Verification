module DP_SOURCE(DP_TL_if tl_if, DP_SINK_if sink_if);















endmodule