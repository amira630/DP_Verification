interface DP_TL_if(clk);
    // ... rest of the code
endinterface