module dp_source(DP_TL_if.DUT tl_if, DP_SINK_if.DUT sink_if);

endmodule
