interface dp_tl_if(input clk);
    string name_1, name_2, name_3;

    // modport DUT (
    //     input clk, reset, valid_in, cin, a, b,
    //     output valid_out, carry, zero, alu
    // );

    
endinterface
