//=======================================================================
// Module: RPTR_EMPTY
// Author: Mohammed Tersawy
// Description: 
// This module implements the read pointer and empty flag logic for an 
// asynchronous FIFO. It includes functionality for gray-to-binary 
// conversion of the write pointer, binary-to-gray conversion of the 
// read pointer, and calculation of the empty flag based on the 
// difference between the read and write pointers. The module ensures 
// proper synchronization between the read and write domains and 
// provides an almost empty signal to indicate when the FIFO is nearly 
// empty. The read address is derived from the binary read pointer, 
// and the empty flag is updated based on the almost empty condition.
//======================================================================

`default_nettype none  // Disable implicit net declarations to avoid unintended wire declarations.

module RPTR_EMPTY 
#( 
   parameter WPTR_WIDTH = 4 , 
   parameter RPTR_WIDTH = 4 , 
   parameter ADDR_WIDTH = 3
)
(
	input  wire                  rinc ,        // Read increment signal to indicate a read operation.
	input  wire [RPTR_WIDTH-1:0] gray_wr_ptr , // Gray-coded write pointer from the write domain.
	input  wire                  rclk ,        // Read clock signal.
	input  wire                  rrst_n ,      // Active-low reset signal for the read domain.
	output wire                  rempty ,      // Empty flag indicating if the FIFO is alnmost empty.
	output wire [ADDR_WIDTH-1:0] r_addr ,      // Read address derived from the binary read pointer.
	output reg  [WPTR_WIDTH-1:0] gray_rd_ptr   // Gray-coded read pointer for synchronization with the write domain.
);

reg [RPTR_WIDTH-1:0] bn_rptr ;      // Binary read pointer.
reg [WPTR_WIDTH-1:0] bn_wptr ;      // Binary write pointer (converted from gray_wr_ptr).
wire                 almost_empty ; // Flag asserted when the FIFO has less than 2 valid data slots.
//reg                 almost_empty ; // Flag asserted when the FIFO has less than 2 valid data slots.
//======================================================================
// SECTION 1: Gray to Binary Conversion for Write Pointer
//======================================================================
always@(posedge rclk or negedge rrst_n) begin
	if(~rrst_n)
	begin
      bn_wptr <= 'b000000;
	end
	else
	begin

    bn_wptr <= {gray_wr_ptr[WPTR_WIDTH-1], 
			    gray_wr_ptr[WPTR_WIDTH-1]^gray_wr_ptr[WPTR_WIDTH-2], 
			    gray_wr_ptr[WPTR_WIDTH-1]^gray_wr_ptr[WPTR_WIDTH-2]^gray_wr_ptr[WPTR_WIDTH-3], 
			    gray_wr_ptr[WPTR_WIDTH-1]^gray_wr_ptr[WPTR_WIDTH-2]^gray_wr_ptr[WPTR_WIDTH-3]^gray_wr_ptr[WPTR_WIDTH-4], 
			    gray_wr_ptr[WPTR_WIDTH-1]^gray_wr_ptr[WPTR_WIDTH-2]^gray_wr_ptr[WPTR_WIDTH-3]^gray_wr_ptr[WPTR_WIDTH-4]^gray_wr_ptr[WPTR_WIDTH-5], 
			    gray_wr_ptr[WPTR_WIDTH-1]^gray_wr_ptr[WPTR_WIDTH-2]^gray_wr_ptr[WPTR_WIDTH-3]^gray_wr_ptr[WPTR_WIDTH-4]^gray_wr_ptr[WPTR_WIDTH-5]^gray_wr_ptr[WPTR_WIDTH-6], 
			    gray_wr_ptr[WPTR_WIDTH-1]^gray_wr_ptr[WPTR_WIDTH-2]^gray_wr_ptr[WPTR_WIDTH-3]^gray_wr_ptr[WPTR_WIDTH-4]^gray_wr_ptr[WPTR_WIDTH-5]^gray_wr_ptr[WPTR_WIDTH-6]^gray_wr_ptr[WPTR_WIDTH-7], 
	     		gray_wr_ptr[WPTR_WIDTH-1]^gray_wr_ptr[WPTR_WIDTH-2]^gray_wr_ptr[WPTR_WIDTH-3]^gray_wr_ptr[WPTR_WIDTH-4]^gray_wr_ptr[WPTR_WIDTH-5]^gray_wr_ptr[WPTR_WIDTH-6]^gray_wr_ptr[WPTR_WIDTH-7]^gray_wr_ptr[WPTR_WIDTH-8], 
		    	gray_wr_ptr[WPTR_WIDTH-1]^gray_wr_ptr[WPTR_WIDTH-2]^gray_wr_ptr[WPTR_WIDTH-3]^gray_wr_ptr[WPTR_WIDTH-4]^gray_wr_ptr[WPTR_WIDTH-5]^gray_wr_ptr[WPTR_WIDTH-6]^gray_wr_ptr[WPTR_WIDTH-7]^gray_wr_ptr[WPTR_WIDTH-8]^gray_wr_ptr[WPTR_WIDTH-9]};
/*
case (gray_wr_ptr)
9'b000000000: bn_wptr <= 9'b000000000;
9'b000000001: bn_wptr <= 9'b000000001;
9'b000000010: bn_wptr <= 9'b000000011;
9'b000000011: bn_wptr <= 9'b000000010;
9'b000000100: bn_wptr <= 9'b000000110;
9'b000000101: bn_wptr <= 9'b000000111;
9'b000000110: bn_wptr <= 9'b000000101;
9'b000000111: bn_wptr <= 9'b000000100;
9'b000001000: bn_wptr <= 9'b000001100;
9'b000001001: bn_wptr <= 9'b000001101;
9'b000001010: bn_wptr <= 9'b000001111;
9'b000001011: bn_wptr <= 9'b000001110;
9'b000001100: bn_wptr <= 9'b000001010;
9'b000001101: bn_wptr <= 9'b000001011;
9'b000001110: bn_wptr <= 9'b000001001;
9'b000001111: bn_wptr <= 9'b000001000;
9'b000010000: bn_wptr <= 9'b000011000;
9'b000010001: bn_wptr <= 9'b000011001;
9'b000010010: bn_wptr <= 9'b000011011;
9'b000010011: bn_wptr <= 9'b000011010;
9'b000010100: bn_wptr <= 9'b000011110;
9'b000010101: bn_wptr <= 9'b000011111;
9'b000010110: bn_wptr <= 9'b000011101;
9'b000010111: bn_wptr <= 9'b000011100;
9'b000011000: bn_wptr <= 9'b000010100;
9'b000011001: bn_wptr <= 9'b000010101;
9'b000011010: bn_wptr <= 9'b000010111;
9'b000011011: bn_wptr <= 9'b000010110;
9'b000011100: bn_wptr <= 9'b000010010;
9'b000011101: bn_wptr <= 9'b000010011;
9'b000011110: bn_wptr <= 9'b000010001;
9'b000011111: bn_wptr <= 9'b000010000;
9'b000100000: bn_wptr <= 9'b000110000;
9'b000100001: bn_wptr <= 9'b000110001;
9'b000100010: bn_wptr <= 9'b000110011;
9'b000100011: bn_wptr <= 9'b000110010;
9'b000100100: bn_wptr <= 9'b000110110;
9'b000100101: bn_wptr <= 9'b000110111;
9'b000100110: bn_wptr <= 9'b000110101;
9'b000100111: bn_wptr <= 9'b000110100;
9'b000101000: bn_wptr <= 9'b000111100;
9'b000101001: bn_wptr <= 9'b000111101;
9'b000101010: bn_wptr <= 9'b000111111;
9'b000101011: bn_wptr <= 9'b000111110;
9'b000101100: bn_wptr <= 9'b000111010;
9'b000101101: bn_wptr <= 9'b000111011;
9'b000101110: bn_wptr <= 9'b000111001;
9'b000101111: bn_wptr <= 9'b000111000;
9'b000110000: bn_wptr <= 9'b000101000;
9'b000110001: bn_wptr <= 9'b000101001;
9'b000110010: bn_wptr <= 9'b000101011;
9'b000110011: bn_wptr <= 9'b000101010;
9'b000110100: bn_wptr <= 9'b000101110;
9'b000110101: bn_wptr <= 9'b000101111;
9'b000110110: bn_wptr <= 9'b000101101;
9'b000110111: bn_wptr <= 9'b000101100;
9'b000111000: bn_wptr <= 9'b000100100;
9'b000111001: bn_wptr <= 9'b000100101;
9'b000111010: bn_wptr <= 9'b000100111;
9'b000111011: bn_wptr <= 9'b000100110;
9'b000111100: bn_wptr <= 9'b000100010;
9'b000111101: bn_wptr <= 9'b000100011;
9'b000111110: bn_wptr <= 9'b000100001;
9'b000111111: bn_wptr <= 9'b000100000;
9'b001000000: bn_wptr <= 9'b001100000;
9'b001000001: bn_wptr <= 9'b001100001;
9'b001000010: bn_wptr <= 9'b001100011;
9'b001000011: bn_wptr <= 9'b001100010;
9'b001000100: bn_wptr <= 9'b001100110;
9'b001000101: bn_wptr <= 9'b001100111;
9'b001000110: bn_wptr <= 9'b001100101;
9'b001000111: bn_wptr <= 9'b001100100;
9'b001001000: bn_wptr <= 9'b001101100;
9'b001001001: bn_wptr <= 9'b001101101;
9'b001001010: bn_wptr <= 9'b001101111;
9'b001001011: bn_wptr <= 9'b001101110;
9'b001001100: bn_wptr <= 9'b001101010;
9'b001001101: bn_wptr <= 9'b001101011;
9'b001001110: bn_wptr <= 9'b001101001;
9'b001001111: bn_wptr <= 9'b001101000;
9'b001010000: bn_wptr <= 9'b001111000;
9'b001010001: bn_wptr <= 9'b001111001;
9'b001010010: bn_wptr <= 9'b001111011;
9'b001010011: bn_wptr <= 9'b001111010;
9'b001010100: bn_wptr <= 9'b001111110;
9'b001010101: bn_wptr <= 9'b001111111;
9'b001010110: bn_wptr <= 9'b001111101;
9'b001010111: bn_wptr <= 9'b001111100;
9'b001011000: bn_wptr <= 9'b001110100;
9'b001011001: bn_wptr <= 9'b001110101;
9'b001011010: bn_wptr <= 9'b001110111;
9'b001011011: bn_wptr <= 9'b001110110;
9'b001011100: bn_wptr <= 9'b001110010;
9'b001011101: bn_wptr <= 9'b001110011;
9'b001011110: bn_wptr <= 9'b001110001;
9'b001011111: bn_wptr <= 9'b001110000;
9'b001100000: bn_wptr <= 9'b001010000;
9'b001100001: bn_wptr <= 9'b001010001;
9'b001100010: bn_wptr <= 9'b001010011;
9'b001100011: bn_wptr <= 9'b001010010;
9'b001100100: bn_wptr <= 9'b001010110;
9'b001100101: bn_wptr <= 9'b001010111;
9'b001100110: bn_wptr <= 9'b001010101;
9'b001100111: bn_wptr <= 9'b001010100;
9'b001101000: bn_wptr <= 9'b001011100;
9'b001101001: bn_wptr <= 9'b001011101;
9'b001101010: bn_wptr <= 9'b001011111;
9'b001101011: bn_wptr <= 9'b001011110;
9'b001101100: bn_wptr <= 9'b001011010;
9'b001101101: bn_wptr <= 9'b001011011;
9'b001101110: bn_wptr <= 9'b001011001;
9'b001101111: bn_wptr <= 9'b001011000;
9'b001110000: bn_wptr <= 9'b001001000;
9'b001110001: bn_wptr <= 9'b001001001;
9'b001110010: bn_wptr <= 9'b001001011;
9'b001110011: bn_wptr <= 9'b001001010;
9'b001110100: bn_wptr <= 9'b001001110;
9'b001110101: bn_wptr <= 9'b001001111;
9'b001110110: bn_wptr <= 9'b001001101;
9'b001110111: bn_wptr <= 9'b001001100;
9'b001111000: bn_wptr <= 9'b001000100;
9'b001111001: bn_wptr <= 9'b001000101;
9'b001111010: bn_wptr <= 9'b001000111;
9'b001111011: bn_wptr <= 9'b001000110;
9'b001111100: bn_wptr <= 9'b001000010;
9'b001111101: bn_wptr <= 9'b001000011;
9'b001111110: bn_wptr <= 9'b001000001;
9'b001111111: bn_wptr <= 9'b001000000;
9'b010000000: bn_wptr <= 9'b011000000;
9'b010000001: bn_wptr <= 9'b011000001;
9'b010000010: bn_wptr <= 9'b011000011;
9'b010000011: bn_wptr <= 9'b011000010;
9'b010000100: bn_wptr <= 9'b011000110;
9'b010000101: bn_wptr <= 9'b011000111;
9'b010000110: bn_wptr <= 9'b011000101;
9'b010000111: bn_wptr <= 9'b011000100;
9'b010001000: bn_wptr <= 9'b011001100;
9'b010001001: bn_wptr <= 9'b011001101;
9'b010001010: bn_wptr <= 9'b011001111;
9'b010001011: bn_wptr <= 9'b011001110;
9'b010001100: bn_wptr <= 9'b011001010;
9'b010001101: bn_wptr <= 9'b011001011;
9'b010001110: bn_wptr <= 9'b011001001;
9'b010001111: bn_wptr <= 9'b011001000;
9'b010010000: bn_wptr <= 9'b011011000;
9'b010010001: bn_wptr <= 9'b011011001;
9'b010010010: bn_wptr <= 9'b011011011;
9'b010010011: bn_wptr <= 9'b011011010;
9'b010010100: bn_wptr <= 9'b011011110;
9'b010010101: bn_wptr <= 9'b011011111;
9'b010010110: bn_wptr <= 9'b011011101;
9'b010010111: bn_wptr <= 9'b011011100;
9'b010011000: bn_wptr <= 9'b011010100;
9'b010011001: bn_wptr <= 9'b011010101;
9'b010011010: bn_wptr <= 9'b011010111;
9'b010011011: bn_wptr <= 9'b011010110;
9'b010011100: bn_wptr <= 9'b011010010;
9'b010011101: bn_wptr <= 9'b011010011;
9'b010011110: bn_wptr <= 9'b011010001;
9'b010011111: bn_wptr <= 9'b011010000;
9'b010100000: bn_wptr <= 9'b011110000;
9'b010100001: bn_wptr <= 9'b011110001;
9'b010100010: bn_wptr <= 9'b011110011;
9'b010100011: bn_wptr <= 9'b011110010;
9'b010100100: bn_wptr <= 9'b011110110;
9'b010100101: bn_wptr <= 9'b011110111;
9'b010100110: bn_wptr <= 9'b011110101;
9'b010100111: bn_wptr <= 9'b011110100;
9'b010101000: bn_wptr <= 9'b011111100;
9'b010101001: bn_wptr <= 9'b011111101;
9'b010101010: bn_wptr <= 9'b011111111;
9'b010101011: bn_wptr <= 9'b011111110;
9'b010101100: bn_wptr <= 9'b011111010;
9'b010101101: bn_wptr <= 9'b011111011;
9'b010101110: bn_wptr <= 9'b011111001;
9'b010101111: bn_wptr <= 9'b011111000;
9'b010110000: bn_wptr <= 9'b011101000;
9'b010110001: bn_wptr <= 9'b011101001;
9'b010110010: bn_wptr <= 9'b011101011;
9'b010110011: bn_wptr <= 9'b011101010;
9'b010110100: bn_wptr <= 9'b011101110;
9'b010110101: bn_wptr <= 9'b011101111;
9'b010110110: bn_wptr <= 9'b011101101;
9'b010110111: bn_wptr <= 9'b011101100;
9'b010111000: bn_wptr <= 9'b011100100;
9'b010111001: bn_wptr <= 9'b011100101;
9'b010111010: bn_wptr <= 9'b011100111;
9'b010111011: bn_wptr <= 9'b011100110;
9'b010111100: bn_wptr <= 9'b011100010;
9'b010111101: bn_wptr <= 9'b011100011;
9'b010111110: bn_wptr <= 9'b011100001;
9'b010111111: bn_wptr <= 9'b011100000;
9'b011000000: bn_wptr <= 9'b010100000;
9'b011000001: bn_wptr <= 9'b010100001;
9'b011000010: bn_wptr <= 9'b010100011;
9'b011000011: bn_wptr <= 9'b010100010;
9'b011000100: bn_wptr <= 9'b010100110;
9'b011000101: bn_wptr <= 9'b010100111;
9'b011000110: bn_wptr <= 9'b010100101;
9'b011000111: bn_wptr <= 9'b010100100;
9'b011001000: bn_wptr <= 9'b010101100;
9'b011001001: bn_wptr <= 9'b010101101;
9'b011001010: bn_wptr <= 9'b010101111;
9'b011001011: bn_wptr <= 9'b010101110;
9'b011001100: bn_wptr <= 9'b010101010;
9'b011001101: bn_wptr <= 9'b010101011;
9'b011001110: bn_wptr <= 9'b010101001;
9'b011001111: bn_wptr <= 9'b010101000;
9'b011010000: bn_wptr <= 9'b010111000;
9'b011010001: bn_wptr <= 9'b010111001;
9'b011010010: bn_wptr <= 9'b010111011;
9'b011010011: bn_wptr <= 9'b010111010;
9'b011010100: bn_wptr <= 9'b010111110;
9'b011010101: bn_wptr <= 9'b010111111;
9'b011010110: bn_wptr <= 9'b010111101;
9'b011010111: bn_wptr <= 9'b010111100;
9'b011011000: bn_wptr <= 9'b010110100;
9'b011011001: bn_wptr <= 9'b010110101;
9'b011011010: bn_wptr <= 9'b010110111;
9'b011011011: bn_wptr <= 9'b010110110;
9'b011011100: bn_wptr <= 9'b010110010;
9'b011011101: bn_wptr <= 9'b010110011;
9'b011011110: bn_wptr <= 9'b010110001;
9'b011011111: bn_wptr <= 9'b010110000;
9'b011100000: bn_wptr <= 9'b010010000;
9'b011100001: bn_wptr <= 9'b010010001;
9'b011100010: bn_wptr <= 9'b010010011;
9'b011100011: bn_wptr <= 9'b010010010;
9'b011100100: bn_wptr <= 9'b010010110;
9'b011100101: bn_wptr <= 9'b010010111;
9'b011100110: bn_wptr <= 9'b010010101;
9'b011100111: bn_wptr <= 9'b010010100;
9'b011101000: bn_wptr <= 9'b010011100;
9'b011101001: bn_wptr <= 9'b010011101;
9'b011101010: bn_wptr <= 9'b010011111;
9'b011101011: bn_wptr <= 9'b010011110;
9'b011101100: bn_wptr <= 9'b010011010;
9'b011101101: bn_wptr <= 9'b010011011;
9'b011101110: bn_wptr <= 9'b010011001;
9'b011101111: bn_wptr <= 9'b010011000;
9'b011110000: bn_wptr <= 9'b010001000;
9'b011110001: bn_wptr <= 9'b010001001;
9'b011110010: bn_wptr <= 9'b010001011;
9'b011110011: bn_wptr <= 9'b010001010;
9'b011110100: bn_wptr <= 9'b010001110;
9'b011110101: bn_wptr <= 9'b010001111;
9'b011110110: bn_wptr <= 9'b010001101;
9'b011110111: bn_wptr <= 9'b010001100;
9'b011111000: bn_wptr <= 9'b010000100;
9'b011111001: bn_wptr <= 9'b010000101;
9'b011111010: bn_wptr <= 9'b010000111;
9'b011111011: bn_wptr <= 9'b010000110;
9'b011111100: bn_wptr <= 9'b010000010;
9'b011111101: bn_wptr <= 9'b010000011;
9'b011111110: bn_wptr <= 9'b010000001;
9'b011111111: bn_wptr <= 9'b010000000;
9'b100000000: bn_wptr <= 9'b110000000;
9'b100000001: bn_wptr <= 9'b110000001;
9'b100000010: bn_wptr <= 9'b110000011;
9'b100000011: bn_wptr <= 9'b110000010;
9'b100000100: bn_wptr <= 9'b110000110;
9'b100000101: bn_wptr <= 9'b110000111;
9'b100000110: bn_wptr <= 9'b110000101;
9'b100000111: bn_wptr <= 9'b110000100;
9'b100001000: bn_wptr <= 9'b110001100;
9'b100001001: bn_wptr <= 9'b110001101;
9'b100001010: bn_wptr <= 9'b110001111;
9'b100001011: bn_wptr <= 9'b110001110;
9'b100001100: bn_wptr <= 9'b110001010;
9'b100001101: bn_wptr <= 9'b110001011;
9'b100001110: bn_wptr <= 9'b110001001;
9'b100001111: bn_wptr <= 9'b110001000;
9'b100010000: bn_wptr <= 9'b110011000;
9'b100010001: bn_wptr <= 9'b110011001;
9'b100010010: bn_wptr <= 9'b110011011;
9'b100010011: bn_wptr <= 9'b110011010;
9'b100010100: bn_wptr <= 9'b110011110;
9'b100010101: bn_wptr <= 9'b110011111;
9'b100010110: bn_wptr <= 9'b110011101;
9'b100010111: bn_wptr <= 9'b110011100;
9'b100011000: bn_wptr <= 9'b110010100;
9'b100011001: bn_wptr <= 9'b110010101;
9'b100011010: bn_wptr <= 9'b110010111;
9'b100011011: bn_wptr <= 9'b110010110;
9'b100011100: bn_wptr <= 9'b110010010;
9'b100011101: bn_wptr <= 9'b110010011;
9'b100011110: bn_wptr <= 9'b110010001;
9'b100011111: bn_wptr <= 9'b110010000;
9'b100100000: bn_wptr <= 9'b110110000;
9'b100100001: bn_wptr <= 9'b110110001;
9'b100100010: bn_wptr <= 9'b110110011;
9'b100100011: bn_wptr <= 9'b110110010;
9'b100100100: bn_wptr <= 9'b110110110;
9'b100100101: bn_wptr <= 9'b110110111;
9'b100100110: bn_wptr <= 9'b110110101;
9'b100100111: bn_wptr <= 9'b110110100;
9'b100101000: bn_wptr <= 9'b110111100;
9'b100101001: bn_wptr <= 9'b110111101;
9'b100101010: bn_wptr <= 9'b110111111;
9'b100101011: bn_wptr <= 9'b110111110;
9'b100101100: bn_wptr <= 9'b110111010;
9'b100101101: bn_wptr <= 9'b110111011;
9'b100101110: bn_wptr <= 9'b110111001;
9'b100101111: bn_wptr <= 9'b110111000;
9'b100110000: bn_wptr <= 9'b110101000;
9'b100110001: bn_wptr <= 9'b110101001;
9'b100110010: bn_wptr <= 9'b110101011;
9'b100110011: bn_wptr <= 9'b110101010;
9'b100110100: bn_wptr <= 9'b110101110;
9'b100110101: bn_wptr <= 9'b110101111;
9'b100110110: bn_wptr <= 9'b110101101;
9'b100110111: bn_wptr <= 9'b110101100;
9'b100111000: bn_wptr <= 9'b110100100;
9'b100111001: bn_wptr <= 9'b110100101;
9'b100111010: bn_wptr <= 9'b110100111;
9'b100111011: bn_wptr <= 9'b110100110;
9'b100111100: bn_wptr <= 9'b110100010;
9'b100111101: bn_wptr <= 9'b110100011;
9'b100111110: bn_wptr <= 9'b110100001;
9'b100111111: bn_wptr <= 9'b110100000;
9'b101000000: bn_wptr <= 9'b111100000;
9'b101000001: bn_wptr <= 9'b111100001;
9'b101000010: bn_wptr <= 9'b111100011;
9'b101000011: bn_wptr <= 9'b111100010;
9'b101000100: bn_wptr <= 9'b111100110;
9'b101000101: bn_wptr <= 9'b111100111;
9'b101000110: bn_wptr <= 9'b111100101;
9'b101000111: bn_wptr <= 9'b111100100;
9'b101001000: bn_wptr <= 9'b111101100;
9'b101001001: bn_wptr <= 9'b111101101;
9'b101001010: bn_wptr <= 9'b111101111;
9'b101001011: bn_wptr <= 9'b111101110;
9'b101001100: bn_wptr <= 9'b111101010;
9'b101001101: bn_wptr <= 9'b111101011;
9'b101001110: bn_wptr <= 9'b111101001;
9'b101001111: bn_wptr <= 9'b111101000;
9'b101010000: bn_wptr <= 9'b111111000;
9'b101010001: bn_wptr <= 9'b111111001;
9'b101010010: bn_wptr <= 9'b111111011;
9'b101010011: bn_wptr <= 9'b111111010;
9'b101010100: bn_wptr <= 9'b111111110;
9'b101010101: bn_wptr <= 9'b111111111;
9'b101010110: bn_wptr <= 9'b111111101;
9'b101010111: bn_wptr <= 9'b111111100;
9'b101011000: bn_wptr <= 9'b111110100;
9'b101011001: bn_wptr <= 9'b111110101;
9'b101011010: bn_wptr <= 9'b111110111;
9'b101011011: bn_wptr <= 9'b111110110;
9'b101011100: bn_wptr <= 9'b111110010;
9'b101011101: bn_wptr <= 9'b111110011;
9'b101011110: bn_wptr <= 9'b111110001;
9'b101011111: bn_wptr <= 9'b111110000;
9'b101100000: bn_wptr <= 9'b111010000;
9'b101100001: bn_wptr <= 9'b111010001;
9'b101100010: bn_wptr <= 9'b111010011;
9'b101100011: bn_wptr <= 9'b111010010;
9'b101100100: bn_wptr <= 9'b111010110;
9'b101100101: bn_wptr <= 9'b111010111;
9'b101100110: bn_wptr <= 9'b111010101;
9'b101100111: bn_wptr <= 9'b111010100;
9'b101101000: bn_wptr <= 9'b111011100;
9'b101101001: bn_wptr <= 9'b111011101;
9'b101101010: bn_wptr <= 9'b111011111;
9'b101101011: bn_wptr <= 9'b111011110;
9'b101101100: bn_wptr <= 9'b111011010;
9'b101101101: bn_wptr <= 9'b111011011;
9'b101101110: bn_wptr <= 9'b111011001;
9'b101101111: bn_wptr <= 9'b111011000;
9'b101110000: bn_wptr <= 9'b111001000;
9'b101110001: bn_wptr <= 9'b111001001;
9'b101110010: bn_wptr <= 9'b111001011;
9'b101110011: bn_wptr <= 9'b111001010;
9'b101110100: bn_wptr <= 9'b111001110;
9'b101110101: bn_wptr <= 9'b111001111;
9'b101110110: bn_wptr <= 9'b111001101;
9'b101110111: bn_wptr <= 9'b111001100;
9'b101111000: bn_wptr <= 9'b111000100;
9'b101111001: bn_wptr <= 9'b111000101;
9'b101111010: bn_wptr <= 9'b111000111;
9'b101111011: bn_wptr <= 9'b111000110;
9'b101111100: bn_wptr <= 9'b111000010;
9'b101111101: bn_wptr <= 9'b111000011;
9'b101111110: bn_wptr <= 9'b111000001;
9'b101111111: bn_wptr <= 9'b111000000;
9'b110000000: bn_wptr <= 9'b101000000;
9'b110000001: bn_wptr <= 9'b101000001;
9'b110000010: bn_wptr <= 9'b101000011;
9'b110000011: bn_wptr <= 9'b101000010;
9'b110000100: bn_wptr <= 9'b101000110;
9'b110000101: bn_wptr <= 9'b101000111;
9'b110000110: bn_wptr <= 9'b101000101;
9'b110000111: bn_wptr <= 9'b101000100;
9'b110001000: bn_wptr <= 9'b101001100;
9'b110001001: bn_wptr <= 9'b101001101;
9'b110001010: bn_wptr <= 9'b101001111;
9'b110001011: bn_wptr <= 9'b101001110;
9'b110001100: bn_wptr <= 9'b101001010;
9'b110001101: bn_wptr <= 9'b101001011;
9'b110001110: bn_wptr <= 9'b101001001;
9'b110001111: bn_wptr <= 9'b101001000;
9'b110010000: bn_wptr <= 9'b101011000;
9'b110010001: bn_wptr <= 9'b101011001;
9'b110010010: bn_wptr <= 9'b101011011;
9'b110010011: bn_wptr <= 9'b101011010;
9'b110010100: bn_wptr <= 9'b101011110;
9'b110010101: bn_wptr <= 9'b101011111;
9'b110010110: bn_wptr <= 9'b101011101;
9'b110010111: bn_wptr <= 9'b101011100;
9'b110011000: bn_wptr <= 9'b101010100;
9'b110011001: bn_wptr <= 9'b101010101;
9'b110011010: bn_wptr <= 9'b101010111;
9'b110011011: bn_wptr <= 9'b101010110;
9'b110011100: bn_wptr <= 9'b101010010;
9'b110011101: bn_wptr <= 9'b101010011;
9'b110011110: bn_wptr <= 9'b101010001;
9'b110011111: bn_wptr <= 9'b101010000;
9'b110100000: bn_wptr <= 9'b101110000;
9'b110100001: bn_wptr <= 9'b101110001;
9'b110100010: bn_wptr <= 9'b101110011;
9'b110100011: bn_wptr <= 9'b101110010;
9'b110100100: bn_wptr <= 9'b101110110;
9'b110100101: bn_wptr <= 9'b101110111;
9'b110100110: bn_wptr <= 9'b101110101;
9'b110100111: bn_wptr <= 9'b101110100;
9'b110101000: bn_wptr <= 9'b101111100;
9'b110101001: bn_wptr <= 9'b101111101;
9'b110101010: bn_wptr <= 9'b101111111;
9'b110101011: bn_wptr <= 9'b101111110;
9'b110101100: bn_wptr <= 9'b101111010;
9'b110101101: bn_wptr <= 9'b101111011;
9'b110101110: bn_wptr <= 9'b101111001;
9'b110101111: bn_wptr <= 9'b101111000;
9'b110110000: bn_wptr <= 9'b101101000;
9'b110110001: bn_wptr <= 9'b101101001;
9'b110110010: bn_wptr <= 9'b101101011;
9'b110110011: bn_wptr <= 9'b101101010;
9'b110110100: bn_wptr <= 9'b101101110;
9'b110110101: bn_wptr <= 9'b101101111;
9'b110110110: bn_wptr <= 9'b101101101;
9'b110110111: bn_wptr <= 9'b101101100;
9'b110111000: bn_wptr <= 9'b101100100;
9'b110111001: bn_wptr <= 9'b101100101;
9'b110111010: bn_wptr <= 9'b101100111;
9'b110111011: bn_wptr <= 9'b101100110;
9'b110111100: bn_wptr <= 9'b101100010;
9'b110111101: bn_wptr <= 9'b101100011;
9'b110111110: bn_wptr <= 9'b101100001;
9'b110111111: bn_wptr <= 9'b101100000;
9'b111000000: bn_wptr <= 9'b100100000;
9'b111000001: bn_wptr <= 9'b100100001;
9'b111000010: bn_wptr <= 9'b100100011;
9'b111000011: bn_wptr <= 9'b100100010;
9'b111000100: bn_wptr <= 9'b100100110;
9'b111000101: bn_wptr <= 9'b100100111;
9'b111000110: bn_wptr <= 9'b100100101;
9'b111000111: bn_wptr <= 9'b100100100;
9'b111001000: bn_wptr <= 9'b100101100;
9'b111001001: bn_wptr <= 9'b100101101;
9'b111001010: bn_wptr <= 9'b100101111;
9'b111001011: bn_wptr <= 9'b100101110;
9'b111001100: bn_wptr <= 9'b100101010;
9'b111001101: bn_wptr <= 9'b100101011;
9'b111001110: bn_wptr <= 9'b100101001;
9'b111001111: bn_wptr <= 9'b100101000;
9'b111010000: bn_wptr <= 9'b100111000;
9'b111010001: bn_wptr <= 9'b100111001;
9'b111010010: bn_wptr <= 9'b100111011;
9'b111010011: bn_wptr <= 9'b100111010;
9'b111010100: bn_wptr <= 9'b100111110;
9'b111010101: bn_wptr <= 9'b100111111;
9'b111010110: bn_wptr <= 9'b100111101;
9'b111010111: bn_wptr <= 9'b100111100;
9'b111011000: bn_wptr <= 9'b100110100;
9'b111011001: bn_wptr <= 9'b100110101;
9'b111011010: bn_wptr <= 9'b100110111;
9'b111011011: bn_wptr <= 9'b100110110;
9'b111011100: bn_wptr <= 9'b100110010;
9'b111011101: bn_wptr <= 9'b100110011;
9'b111011110: bn_wptr <= 9'b100110001;
9'b111011111: bn_wptr <= 9'b100110000;
9'b111100000: bn_wptr <= 9'b100010000;
9'b111100001: bn_wptr <= 9'b100010001;
9'b111100010: bn_wptr <= 9'b100010011;
9'b111100011: bn_wptr <= 9'b100010010;
9'b111100100: bn_wptr <= 9'b100010110;
9'b111100101: bn_wptr <= 9'b100010111;
9'b111100110: bn_wptr <= 9'b100010101;
9'b111100111: bn_wptr <= 9'b100010100;
9'b111101000: bn_wptr <= 9'b100011100;
9'b111101001: bn_wptr <= 9'b100011101;
9'b111101010: bn_wptr <= 9'b100011111;
9'b111101011: bn_wptr <= 9'b100011110;
9'b111101100: bn_wptr <= 9'b100011010;
9'b111101101: bn_wptr <= 9'b100011011;
9'b111101110: bn_wptr <= 9'b100011001;
9'b111101111: bn_wptr <= 9'b100011000;
9'b111110000: bn_wptr <= 9'b100001000;
9'b111110001: bn_wptr <= 9'b100001001;
9'b111110010: bn_wptr <= 9'b100001011;
9'b111110011: bn_wptr <= 9'b100001010;
9'b111110100: bn_wptr <= 9'b100001110;
9'b111110101: bn_wptr <= 9'b100001111;
9'b111110110: bn_wptr <= 9'b100001101;
9'b111110111: bn_wptr <= 9'b100001100;
9'b111111000: bn_wptr <= 9'b100000100;
9'b111111001: bn_wptr <= 9'b100000101;
9'b111111010: bn_wptr <= 9'b100000111;
9'b111111011: bn_wptr <= 9'b100000110;
9'b111111100: bn_wptr <= 9'b100000010;
9'b111111101: bn_wptr <= 9'b100000011;
9'b111111110: bn_wptr <= 9'b100000001;
9'b111111111: bn_wptr <= 9'b100000000;
endcase
*/

/*			
case (gray_wr_ptr)
8'b0000000: bn_wptr <= 8'b0000000;
8'b0000001: bn_wptr <= 8'b0000001;
8'b0000011: bn_wptr <= 8'b0000010;
8'b0000010: bn_wptr <= 8'b0000011;
8'b0000110: bn_wptr <= 8'b0000100;
8'b0000111: bn_wptr <= 8'b0000101;
8'b0000101: bn_wptr <= 8'b0000110;
8'b0000100: bn_wptr <= 8'b0000111;
8'b0001100: bn_wptr <= 8'b0001000;
8'b0001101: bn_wptr <= 8'b0001001;
8'b0001111: bn_wptr <= 8'b0001010;
8'b0001110: bn_wptr <= 8'b0001011;
8'b0001010: bn_wptr <= 8'b0001100;
8'b0001011: bn_wptr <= 8'b0001101;
8'b0001001: bn_wptr <= 8'b0001110;
8'b0001000: bn_wptr <= 8'b0001111;

8'b0011000: bn_wptr <= 8'b0010000;
8'b0011001: bn_wptr <= 8'b0010001;
8'b0011011: bn_wptr <= 8'b0010010;
8'b0011010: bn_wptr <= 8'b0010011;
8'b0011110: bn_wptr <= 8'b0010100;
8'b0011111: bn_wptr <= 8'b0010101;
8'b0011101: bn_wptr <= 8'b0010110;
8'b0011100: bn_wptr <= 8'b0010111;
8'b0010100: bn_wptr <= 8'b0011000;
8'b0010101: bn_wptr <= 8'b0011001;
8'b0010111: bn_wptr <= 8'b0011010;
8'b0010110: bn_wptr <= 8'b0011011;
8'b0010010: bn_wptr <= 8'b0011100;
8'b0010011: bn_wptr <= 8'b0011101;
8'b0010001: bn_wptr <= 8'b0011110;
8'b0010000: bn_wptr <= 8'b0011111;

8'b0011000: bn_wptr <= 8'b0100000;
8'b0011001: bn_wptr <= 8'b0100001;
8'b0011011: bn_wptr <= 8'b0100010;
8'b0011010: bn_wptr <= 8'b0100011;
8'b0011110: bn_wptr <= 8'b0100100;
8'b0011111: bn_wptr <= 8'b0100101;
8'b0011101: bn_wptr <= 8'b0100110;
8'b0011100: bn_wptr <= 8'b0100111;
8'b0010100: bn_wptr <= 8'b0101000;
8'b0010101: bn_wptr <= 8'b0101001;
8'b0010111: bn_wptr <= 8'b0101010;
8'b0010110: bn_wptr <= 8'b0101011;
8'b0010010: bn_wptr <= 8'b0101100;
8'b0010011: bn_wptr <= 8'b0101101;
8'b0010001: bn_wptr <= 8'b0101110;
8'b0010000: bn_wptr <= 8'b0101111;

8'b0110000: bn_wptr <= 8'b0100000;
8'b0110001: bn_wptr <= 8'b0100001;
8'b0110011: bn_wptr <= 8'b0100010;
8'b0110010: bn_wptr <= 8'b0100011;
8'b0110110: bn_wptr <= 8'b0100100;
8'b0110111: bn_wptr <= 8'b0100101;
8'b0110101: bn_wptr <= 8'b0100110;
8'b0110100: bn_wptr <= 8'b0100111;
8'b0111100: bn_wptr <= 8'b0101000;
8'b0111101: bn_wptr <= 8'b0101001;
8'b0111111: bn_wptr <= 8'b0101010;
8'b0111110: bn_wptr <= 8'b0101011;
8'b0111010: bn_wptr <= 8'b0101100;
8'b0111011: bn_wptr <= 8'b0101101;
8'b0111001: bn_wptr <= 8'b0101110;
8'b0111000: bn_wptr <= 8'b0101111;

8'b1101000: bn_wptr <= 8'b0110000;
8'b1101001: bn_wptr <= 8'b0110001;
8'b1101011: bn_wptr <= 8'b0110010;
8'b1101010: bn_wptr <= 8'b0110011;
8'b1101110: bn_wptr <= 8'b0110100;
8'b1101111: bn_wptr <= 8'b0110101;
8'b1101101: bn_wptr <= 8'b0110110;
8'b1101100: bn_wptr <= 8'b0110111;
8'b1100100: bn_wptr <= 8'b0111000;
8'b1100101: bn_wptr <= 8'b0111001;
8'b1100111: bn_wptr <= 8'b0111010;
8'b1100110: bn_wptr <= 8'b0111011;
8'b1100010: bn_wptr <= 8'b0111100;
8'b1100011: bn_wptr <= 8'b0111101;
8'b1100001: bn_wptr <= 8'b0111110;
8'b1100000: bn_wptr <= 8'b0111111;

8'b1111000: bn_wptr <= 8'b1000000;
8'b1111001: bn_wptr <= 8'b1000001;
8'b1111011: bn_wptr <= 8'b1000010;
8'b1111010: bn_wptr <= 8'b1000011;
8'b1111110: bn_wptr <= 8'b1000100;
8'b1111111: bn_wptr <= 8'b1000101;
8'b1111101: bn_wptr <= 8'b1000110;
8'b1111100: bn_wptr <= 8'b1000111;
8'b1110100: bn_wptr <= 8'b1001000;
8'b1110101: bn_wptr <= 8'b1001001;
8'b1110111: bn_wptr <= 8'b1001010;
8'b1110110: bn_wptr <= 8'b1001011;
8'b1110010: bn_wptr <= 8'b1001100;
8'b1110011: bn_wptr <= 8'b1001101;
8'b1110001: bn_wptr <= 8'b1001110;
8'b1110000: bn_wptr <= 8'b1001111;

8'b1010000: bn_wptr <= 8'b1010000;
8'b1010001: bn_wptr <= 8'b1010001;
8'b1010011: bn_wptr <= 8'b1010010;
8'b1010010: bn_wptr <= 8'b1010011;
8'b1010110: bn_wptr <= 8'b1010100;
8'b1010111: bn_wptr <= 8'b1010101;
8'b1010101: bn_wptr <= 8'b1010110;
8'b1010100: bn_wptr <= 8'b1010111;
8'b1011100: bn_wptr <= 8'b1011000;
8'b1011101: bn_wptr <= 8'b1011001;
8'b1011111: bn_wptr <= 8'b1011010;
8'b1011110: bn_wptr <= 8'b1011011;
8'b1011010: bn_wptr <= 8'b1011100;
8'b1011011: bn_wptr <= 8'b1011101;
8'b1011001: bn_wptr <= 8'b1011110;
8'b1011000: bn_wptr <= 8'b1011111;

8'b1001000: bn_wptr <= 8'b1100000;
8'b1001001: bn_wptr <= 8'b1100001;
8'b1001011: bn_wptr <= 8'b1100010;
8'b1001010: bn_wptr <= 8'b1100011;
8'b1001110: bn_wptr <= 8'b1100100;
8'b1001111: bn_wptr <= 8'b1100101;
8'b1001101: bn_wptr <= 8'b1100110;
8'b1001100: bn_wptr <= 8'b1100111;
8'b1000100: bn_wptr <= 8'b1101000;
8'b1000101: bn_wptr <= 8'b1101001;
8'b1000111: bn_wptr <= 8'b1101010;
8'b1000110: bn_wptr <= 8'b1101011;
8'b1000010: bn_wptr <= 8'b1101100;
8'b1000011: bn_wptr <= 8'b1101101;
8'b1000001: bn_wptr <= 8'b1101110;
8'b1000000: bn_wptr <= 8'b1101111;

8'b0001000: bn_wptr <= 8'b1110000;
8'b0001001: bn_wptr <= 8'b1110001;
8'b0001011: bn_wptr <= 8'b1110010;
8'b0001010: bn_wptr <= 8'b1110011;
8'b0001110: bn_wptr <= 8'b1110100;
8'b0001111: bn_wptr <= 8'b1110101;
8'b0001101: bn_wptr <= 8'b1110110;
8'b0001100: bn_wptr <= 8'b1110111;
8'b0000100: bn_wptr <= 8'b1111000;
8'b0000101: bn_wptr <= 8'b1111001;
8'b0000111: bn_wptr <= 8'b1111010;
8'b0000110: bn_wptr <= 8'b1111011;
8'b0000010: bn_wptr <= 8'b1111100;
8'b0000011: bn_wptr <= 8'b1111101;
8'b0000001: bn_wptr <= 8'b1111110;
8'b0000000: bn_wptr <= 8'b1111111;

// Complete 8-bit bit reversal mapping (256 cases)
// Format: 8'bABCDEFGH maps to 8'bHGFEDCBA

// Cases 0-15
8'b00000000: bn_wptr <= 8'b00000000;
8'b00000001: bn_wptr <= 8'b10000000;
8'b00000010: bn_wptr <= 8'b01000000;
8'b00000011: bn_wptr <= 8'b11000000;
8'b00000100: bn_wptr <= 8'b00100000;
8'b00000101: bn_wptr <= 8'b10100000;
8'b00000110: bn_wptr <= 8'b01100000;
8'b00000111: bn_wptr <= 8'b11100000;
8'b00001000: bn_wptr <= 8'b00010000;
8'b00001001: bn_wptr <= 8'b10010000;
8'b00001010: bn_wptr <= 8'b01010000;
8'b00001011: bn_wptr <= 8'b11010000;
8'b00001100: bn_wptr <= 8'b00110000;
8'b00001101: bn_wptr <= 8'b10110000;
8'b00001110: bn_wptr <= 8'b01110000;
8'b00001111: bn_wptr <= 8'b11110000;

// Cases 16-31
8'b00010000: bn_wptr <= 8'b00001000;
8'b00010001: bn_wptr <= 8'b10001000;
8'b00010010: bn_wptr <= 8'b01001000;
8'b00010011: bn_wptr <= 8'b11001000;
8'b00010100: bn_wptr <= 8'b00101000;
8'b00010101: bn_wptr <= 8'b10101000;
8'b00010110: bn_wptr <= 8'b01101000;
8'b00010111: bn_wptr <= 8'b11101000;
8'b00011000: bn_wptr <= 8'b00011000;
8'b00011001: bn_wptr <= 8'b10011000;
8'b00011010: bn_wptr <= 8'b01011000;
8'b00011011: bn_wptr <= 8'b11011000;
8'b00011100: bn_wptr <= 8'b00111000;
8'b00011101: bn_wptr <= 8'b10111000;
8'b00011110: bn_wptr <= 8'b01111000;
8'b00011111: bn_wptr <= 8'b11111000;

// Cases 32-48
8'b00100000: bn_wptr <= 8'b00000100;
8'b00100001: bn_wptr <= 8'b10000100;
8'b00100010: bn_wptr <= 8'b01000100;
8'b00100011: bn_wptr <= 8'b11000100;
8'b00100100: bn_wptr <= 8'b00100100;
8'b00100101: bn_wptr <= 8'b10100100;
8'b00100110: bn_wptr <= 8'b01100100;
8'b00100111: bn_wptr <= 8'b11100100;
8'b00101000: bn_wptr <= 8'b00010100;
8'b00101001: bn_wptr <= 8'b10010100;
8'b00101010: bn_wptr <= 8'b01010100;
8'b00101011: bn_wptr <= 8'b11010100;
8'b00101100: bn_wptr <= 8'b00110100;
8'b00101101: bn_wptr <= 8'b10110100;
8'b00101110: bn_wptr <= 8'b01110100;
8'b00101111: bn_wptr <= 8'b11110100;

// Cases 48-63
8'b00110000: bn_wptr <= 8'b00001100;
8'b00110001: bn_wptr <= 8'b10001100;
8'b00110010: bn_wptr <= 8'b01001100;
8'b00110011: bn_wptr <= 8'b11001100;
8'b00110100: bn_wptr <= 8'b00101100;
8'b00110101: bn_wptr <= 8'b10101100;
8'b00110110: bn_wptr <= 8'b01101100;
8'b00110111: bn_wptr <= 8'b11101100;
8'b00111000: bn_wptr <= 8'b00011100;
8'b00111001: bn_wptr <= 8'b10011100;
8'b00111010: bn_wptr <= 8'b01011100;
8'b00111011: bn_wptr <= 8'b11011100;
8'b00111100: bn_wptr <= 8'b00111100;
8'b00111101: bn_wptr <= 8'b10111100;
8'b00111110: bn_wptr <= 8'b01111100;
8'b00111111: bn_wptr <= 8'b11111100;

// Cases 64-89
8'b01000000: bn_wptr <= 8'b00000010;
8'b01000001: bn_wptr <= 8'b10000010;
8'b01000010: bn_wptr <= 8'b01000010;
8'b01000011: bn_wptr <= 8'b11000010;
8'b01000100: bn_wptr <= 8'b00100010;
8'b01000101: bn_wptr <= 8'b10100010;
8'b01000110: bn_wptr <= 8'b01100010;
8'b01000111: bn_wptr <= 8'b11100010;
8'b01001000: bn_wptr <= 8'b00010010;
8'b01001001: bn_wptr <= 8'b10010010;
8'b01001010: bn_wptr <= 8'b01010010;
8'b01001011: bn_wptr <= 8'b11010010;
8'b01001100: bn_wptr <= 8'b00110010;
8'b01001101: bn_wptr <= 8'b10110010;
8'b01001110: bn_wptr <= 8'b01110010;
8'b01001111: bn_wptr <= 8'b11110010;

// Cases 80-95
8'b01010000: bn_wptr <= 8'b00001010;
8'b01010001: bn_wptr <= 8'b10001010;
8'b01010010: bn_wptr <= 8'b01001010;
8'b01010011: bn_wptr <= 8'b11001010;
8'b01010100: bn_wptr <= 8'b00101010;
8'b01010101: bn_wptr <= 8'b10101010;
8'b01010110: bn_wptr <= 8'b01101010;
8'b01010111: bn_wptr <= 8'b11101010;
8'b01011000: bn_wptr <= 8'b00011010;
8'b01011001: bn_wptr <= 8'b10011010;
8'b01011010: bn_wptr <= 8'b01011010;
8'b01011011: bn_wptr <= 8'b11011010;
8'b01011100: bn_wptr <= 8'b00111010;
8'b01011101: bn_wptr <= 8'b10111010;
8'b01011110: bn_wptr <= 8'b01111010;
8'b01011111: bn_wptr <= 8'b11111010;

// Cases 96-111
8'b01100000: bn_wptr <= 8'b00000110;
8'b01100001: bn_wptr <= 8'b10000110;
8'b01100010: bn_wptr <= 8'b01000110;
8'b01100011: bn_wptr <= 8'b11000110;
8'b01100100: bn_wptr <= 8'b00100110;
8'b01100101: bn_wptr <= 8'b10100110;
8'b01100110: bn_wptr <= 8'b01100110;
8'b01100111: bn_wptr <= 8'b11100110;
8'b01101000: bn_wptr <= 8'b00010110;
8'b01101001: bn_wptr <= 8'b10010110;
8'b01101010: bn_wptr <= 8'b01010110;
8'b01101011: bn_wptr <= 8'b11010110;
8'b01101100: bn_wptr <= 8'b00110110;
8'b01101101: bn_wptr <= 8'b10110110;
8'b01101110: bn_wptr <= 8'b01110110;
8'b01101111: bn_wptr <= 8'b11110110;

// Cases 112-128
8'b01110000: bn_wptr <= 8'b00001110;
8'b01110001: bn_wptr <= 8'b10001110;
8'b01110010: bn_wptr <= 8'b01001110;
8'b01110011: bn_wptr <= 8'b11001110;
8'b01110100: bn_wptr <= 8'b00101110;
8'b01110101: bn_wptr <= 8'b10101110;
8'b01110110: bn_wptr <= 8'b01101110;
8'b01110111: bn_wptr <= 8'b11101110;
8'b01111000: bn_wptr <= 8'b00011110;
8'b01111001: bn_wptr <= 8'b10011110;
8'b01111010: bn_wptr <= 8'b01011110;
8'b01111011: bn_wptr <= 8'b11011110;
8'b01111100: bn_wptr <= 8'b00111110;
8'b01111101: bn_wptr <= 8'b10111110;
8'b01111110: bn_wptr <= 8'b01111110;
8'b01111111: bn_wptr <= 8'b11111110;

// Cases 128-143
8'b10000000: bn_wptr <= 8'b00000001;
8'b10000001: bn_wptr <= 8'b10000001;
8'b10000010: bn_wptr <= 8'b01000001;
8'b10000011: bn_wptr <= 8'b11000001;
8'b10000100: bn_wptr <= 8'b00100001;
8'b10000101: bn_wptr <= 8'b10100001;
8'b10000110: bn_wptr <= 8'b01100001;
8'b10000111: bn_wptr <= 8'b11100001;
8'b10001000: bn_wptr <= 8'b00010001;
8'b10001001: bn_wptr <= 8'b10010001;
8'b10001010: bn_wptr <= 8'b01010001;
8'b10001011: bn_wptr <= 8'b11010001;
8'b10001100: bn_wptr <= 8'b00110001;
8'b10001101: bn_wptr <= 8'b10110001;
8'b10001110: bn_wptr <= 8'b01110001;
8'b10001111: bn_wptr <= 8'b11110001;

// Cases 144-159
8'b10010000: bn_wptr <= 8'b00001001;
8'b10010001: bn_wptr <= 8'b10001001;
8'b10010010: bn_wptr <= 8'b01001001;
8'b10010011: bn_wptr <= 8'b11001001;
8'b10010100: bn_wptr <= 8'b00101001;
8'b10010101: bn_wptr <= 8'b10101001;
8'b10010110: bn_wptr <= 8'b01101001;
8'b10010111: bn_wptr <= 8'b11101001;
8'b10011000: bn_wptr <= 8'b00011001;
8'b10011001: bn_wptr <= 8'b10011001;
8'b10011010: bn_wptr <= 8'b01011001;
8'b10011011: bn_wptr <= 8'b11011001;
8'b10011100: bn_wptr <= 8'b00111001;
8'b10011101: bn_wptr <= 8'b10111001;
8'b10011110: bn_wptr <= 8'b01111001;
8'b10011111: bn_wptr <= 8'b11111001;

// Cases 160-185
8'b10100000: bn_wptr <= 8'b00000101;
8'b10100001: bn_wptr <= 8'b10000101;
8'b10100010: bn_wptr <= 8'b01000101;
8'b10100011: bn_wptr <= 8'b11000101;
8'b10100100: bn_wptr <= 8'b00100101;
8'b10100101: bn_wptr <= 8'b10100101;
8'b10100110: bn_wptr <= 8'b01100101;
8'b10100111: bn_wptr <= 8'b11100101;
8'b10101000: bn_wptr <= 8'b00010101;
8'b10101001: bn_wptr <= 8'b10010101;
8'b10101010: bn_wptr <= 8'b01010101;
8'b10101011: bn_wptr <= 8'b11010101;
8'b10101100: bn_wptr <= 8'b00110101;
8'b10101101: bn_wptr <= 8'b10110101;
8'b10101110: bn_wptr <= 8'b01110101;
8'b10101111: bn_wptr <= 8'b11110101;

// Cases 186-191
8'b10110000: bn_wptr <= 8'b00001101;
8'b10110001: bn_wptr <= 8'b10001101;
8'b10110010: bn_wptr <= 8'b01001101;
8'b10110011: bn_wptr <= 8'b11001101;
8'b10110100: bn_wptr <= 8'b00101101;
8'b10110101: bn_wptr <= 8'b10101101;
8'b10110110: bn_wptr <= 8'b01101101;
8'b10110111: bn_wptr <= 8'b11101101;
8'b10111000: bn_wptr <= 8'b00011101;
8'b10111001: bn_wptr <= 8'b10011101;
8'b10111010: bn_wptr <= 8'b01011101;
8'b10111011: bn_wptr <= 8'b11011101;
8'b10111100: bn_wptr <= 8'b00111101;
8'b10111101: bn_wptr <= 8'b10111101;
8'b10111110: bn_wptr <= 8'b01111101;
8'b10111111: bn_wptr <= 8'b11111101;

// Cases 192-208
8'b11000000: bn_wptr <= 8'b00000011;
8'b11000001: bn_wptr <= 8'b10000011;
8'b11000010: bn_wptr <= 8'b01000011;
8'b11000011: bn_wptr <= 8'b11000011;
8'b11000100: bn_wptr <= 8'b00100011;
8'b11000101: bn_wptr <= 8'b10100011;
8'b11000110: bn_wptr <= 8'b01100011;
8'b11000111: bn_wptr <= 8'b11100011;
8'b11001000: bn_wptr <= 8'b00010011;
8'b11001001: bn_wptr <= 8'b10010011;
8'b11001010: bn_wptr <= 8'b01010011;
8'b11001011: bn_wptr <= 8'b11010011;
8'b11001100: bn_wptr <= 8'b00110011;
8'b11001101: bn_wptr <= 8'b10110011;
8'b11001110: bn_wptr <= 8'b01110011;
8'b11001111: bn_wptr <= 8'b11110011;

// Cases 208-223
8'b11010000: bn_wptr <= 8'b00001011;
8'b11010001: bn_wptr <= 8'b10001011;
8'b11010010: bn_wptr <= 8'b01001011;
8'b11010011: bn_wptr <= 8'b11001011;
8'b11010100: bn_wptr <= 8'b00101011;
8'b11010101: bn_wptr <= 8'b10101011;
8'b11010110: bn_wptr <= 8'b01101011;
8'b11010111: bn_wptr <= 8'b11101011;
8'b11011000: bn_wptr <= 8'b00011011;
8'b11011001: bn_wptr <= 8'b10011011;
8'b11011010: bn_wptr <= 8'b01011011;
8'b11011011: bn_wptr <= 8'b11011011;
8'b11011100: bn_wptr <= 8'b00111011;
8'b11011101: bn_wptr <= 8'b10111011;
8'b11011110: bn_wptr <= 8'b01111011;
8'b11011111: bn_wptr <= 8'b11111011;

// Cases 224-239
8'b11100000: bn_wptr <= 8'b00000111;
8'b11100001: bn_wptr <= 8'b10000111;
8'b11100010: bn_wptr <= 8'b01000111;
8'b11100011: bn_wptr <= 8'b11000111;
8'b11100100: bn_wptr <= 8'b00100111;
8'b11100101: bn_wptr <= 8'b10100111;
8'b11100110: bn_wptr <= 8'b01100111;
8'b11100111: bn_wptr <= 8'b11100111;
8'b11101000: bn_wptr <= 8'b00010111;
8'b11101001: bn_wptr <= 8'b10010111;
8'b11101010: bn_wptr <= 8'b01010111;
8'b11101011: bn_wptr <= 8'b11010111;
8'b11101100: bn_wptr <= 8'b00110111;
8'b11101101: bn_wptr <= 8'b10110111;
8'b11101110: bn_wptr <= 8'b01110111;
8'b11101111: bn_wptr <= 8'b11110111;

// Cases 240-255
8'b11110000: bn_wptr <= 8'b00001111;
8'b11110001: bn_wptr <= 8'b10001111;
8'b11110010: bn_wptr <= 8'b01001111;
8'b11110011: bn_wptr <= 8'b11001111;
8'b11110100: bn_wptr <= 8'b00101111;
8'b11110101: bn_wptr <= 8'b10101111;
8'b11110110: bn_wptr <= 8'b01101111;
8'b11110111: bn_wptr <= 8'b11101111;
8'b11111000: bn_wptr <= 8'b00011111;
8'b11111001: bn_wptr <= 8'b10011111;
8'b11111010: bn_wptr <= 8'b01011111;
8'b11111011: bn_wptr <= 8'b11011111;
8'b11111100: bn_wptr <= 8'b00111111;
8'b11111101: bn_wptr <= 8'b10111111;
8'b11111110: bn_wptr <= 8'b01111111;
8'b11111111: bn_wptr <= 8'b11111111;
	endcase
	*/
//bn_wptr <= gray_wr_ptr ^ (gray_wr_ptr >> 1);
	end
end


//======================================================================
// SECTION 2: Almost Empty Signal Calculation
//======================================================================
assign almost_empty = ((bn_wptr - bn_rptr) <= 1'd1); // Check if the difference between write and read pointers is less than 2 slots.
assign rempty = almost_empty ; // Set the empty flag based on the almost_empty condition.
/*
always @(posedge rclk or negedge rrst_n) begin 
	// Update the binary read pointer (bn_rptr) on the rising edge of the read clock or reset.
	if(~rrst_n) 
	begin
		almost_empty <= 1'b0 ; // Reset the binary read pointer to 0.
	end 
	else if ( (bn_wptr - bn_rptr) <= 1 ) 
	begin
		almost_empty <= 1'b1 ; // Increment the binary read pointer by 2 if rinc is asserted and FIFO is not almost empty.
	end 
	else
	begin
       almost_empty <= 1'b0 ;
	end

end
*/
//======================================================================
// SECTION 3: Binary Read Pointer Update
//======================================================================
always @(posedge rclk or negedge rrst_n) begin 
	// Update the binary read pointer (bn_rptr) on the rising edge of the read clock or reset.
	if(~rrst_n) 
	begin
		bn_rptr <= 'b0 ; // Reset the binary read pointer to 0.
	end 
	else 
	if ( rinc == 1'b1 && !almost_empty ) 
	begin
		bn_rptr <= bn_rptr + 'd2 ; // Increment the binary read pointer by 2 if rinc is asserted and FIFO is not almost empty.
	end 
end

//======================================================================
// SECTION 4: Read Address Calculation
//======================================================================
assign r_addr = bn_rptr[ADDR_WIDTH-1:0] ; // Extract the read address from the binary read pointer (excluding the MSB).

//======================================================================
// SECTION 5: Gray-Coded Read Pointer Update
//======================================================================
always @(posedge rclk or negedge rrst_n ) begin
	// Update the gray-coded read pointer (gray_rd_ptr) on the rising edge of the read clock or reset.
	if (~rrst_n) 
	begin
		gray_rd_ptr <= 'b0 ; // Reset the gray-coded read pointer to 0.
	end 
	else 
	begin
		gray_rd_ptr <= bn_rptr ^ (bn_rptr >> 1); // Convert the binary read pointer to gray code.
	end
end

endmodule 

`resetall  // Reset all compiler directives to their default values.
