SINK SINK SINK SINK
SINK SINK SINK SINK SINK