package dp_dpcd_reg_pkg;    
    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Any further package imports:
    //import test_parameters_pkg::*;
    import dp_dpcd_reg_file_receiver_capability_pkg::*;

    // Includes:
    `include "dp_dpcd_reg_block.svh"
endpackage