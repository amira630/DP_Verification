package dp_sink_agent_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Includes:
    `include "dp_source_config.svh"
    `include "dp_sink_sequence_item.svh"
    `include "dp_sink_sequencer.svh"
    `include "dp_sink_driver.svh"
    `include "dp_sink_monitor.svh"
    `include "dp_sink_agent.svh"

endpackage
