package dp_transactions_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Any further package imports:
    import test_parameters_pkg::*;
    
    // Includes:
    `include "dp_source_config.svh"
    `include "dp_tl_spm_sequence_item.svh"
    `include "dp_tl_lpm_sequence_item.svh"
    `include "dp_sink_sequence_item.svh"

endpackage