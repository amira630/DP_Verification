package test_parameters_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "test_parameters.svh"
    
endpackage